library verilog;
use verilog.vl_types.all;
entity mux_test_vlg_vec_tst is
end mux_test_vlg_vec_tst;
