library verilog;
use verilog.vl_types.all;
entity FullBaseStation_vlg_vec_tst is
end FullBaseStation_vlg_vec_tst;
